module mux16x1_TB();
    reg [3:0] S;
    reg [15:0] D;
    wire Y;

    mux16x1 uut (.S(S), .D(D), .Y(Y));

    initial begin
        D[15:0] = 16'b0000000000000000;
        
        S = 4'b0000; #10;
        D[0] = 1; #10;
        S = 4'b0001; #10;
        D[1] = 1; #10;
        S = 4'b0010; #10;
        D[2] = 1; #10;
        S = 4'b0011; #10;
        D[3] = 1; #10;
        S = 4'b0100; #10;
        D[4] = 1; #10;
        S = 4'b0101; #10;
        D[5] = 1; #10;
        S = 4'b0110; #10;
        D[6] = 1; #10;
        S = 4'b0111; #10;
        D[7] = 1; #10;
        S = 4'b1000; #10;
        D[8] = 1; #10;
        S = 4'b1001; #10;
        D[9] = 1; #10;
        S = 4'b1010; #10;
        D[10] = 1; #10;
        S = 4'b1011; #10;
        D[11] = 1; #10;
        S = 4'b1100; #10;
        D[12] = 1; #10;
        S = 4'b1101; #10;
        D[13] = 1; #10;
        S = 4'b1110; #10;
        D[14] = 1; #10;
        S = 4'b1111; #10;
        D[15] = 1; #10;

        $stop;
    end

    initial begin
        $monitor("Tempo = %0t | S = %b | Y = %b | D = %b", $time, S, Y, D[15:0]);
    end
endmodule