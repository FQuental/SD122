module priori16_tb ();
    reg [15:0] in;
    wire [3:0] out;

    priori16x4 uut (.in(in), .out(out));
    initial begin
        $monitor("in = %b, out = %b", in , out);
        in = 16'b0000000000000001; #10; // 00 -> 0000
        in = 16'b0000000000000010; #10; // 01 -> 0001
        in = 16'b0000000000000100; #10; // 02 -> 0010
        in = 16'b0000000000001000; #10; // 03 -> 0011
        in = 16'b0000000000010000; #10; // 04 -> 0100
        in = 16'b0000000000100000; #10; // 05 -> 0101
        in = 16'b0000000001000000; #10; // 06 -> 0110
        in = 16'b0000000010000000; #10; // 07 -> 0111
        in = 16'b0000000100000000; #10; // 08 -> 1000
        in = 16'b0000001000000000; #10; // 09 -> 1001
        in = 16'b0000010000000000; #10; // 10 -> 1010
        in = 16'b0000100000000000; #10; // 11 -> 1011
        in = 16'b0001000000000000; #10; // 12 -> 1100
        in = 16'b0010000000000000; #10; // 13 -> 1101
        in = 16'b0100000000000000; #10; // 14 -> 1110
        in = 16'b1000000000000000; #10; // 15 -> 1111
        $stop;
    end
endmodule