module decode4x16_tb_att2 ();
    reg [3:0] in;
    wire [15:0] out;

    code4x16 uut (.in(in), .out(out));
    initial begin
        $monitor("in = %b, out = %b", in , out);
        in = 4'b1111; #10; // 00 -> 0000
        in = 4'b1110; #10; // 01 -> 0001
        in = 4'b1101; #10; // 02 -> 0010
        in = 4'b1100; #10; // 03 -> 0011
        in = 4'b1011; #10; // 04 -> 0100
        in = 4'b1010; #10; // 05 -> 0101
        in = 4'b1001; #10; // 06 -> 0110
        in = 4'b1000; #10; // 07 -> 0111
        in = 4'b0111; #10; // 08 -> 1000
        in = 4'b0110; #10; // 09 -> 1001
        in = 4'b0101; #10; // 10 -> 1010
        in = 4'b0100; #10; // 11 -> 1011
        in = 4'b0011; #10; // 12 -> 1100
        in = 4'b0010; #10; // 13 -> 1101
        in = 4'b0001; #10; // 14 -> 1110
        in = 4'b0000; #10; // 15 -> 1111
        $stop;
    end
endmodule